// Copyright (c) 2024 Ethan Sifferman.
// All rights reserved. Distribution Prohibited.

package muladd_pkg;

typedef enum logic [1:0] {
    IDLE,
    MUL,
    ADD
} state_t;

endpackage
